//top level snes, calls snes decoder
