//decodes ps2 input, encodes it into desired format
