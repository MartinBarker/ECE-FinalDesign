//gets input from ps2 and snes, translates that input to VGA changes. 
//creates vga display simulation (?)
