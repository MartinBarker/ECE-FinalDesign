//decodes snes input and translates it to desired format
