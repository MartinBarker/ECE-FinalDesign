//top level ps2 , calls ps2 decoder file.
//gets input from ps2 controller, translates input into readable form (or
//number?)
