//brings everything together in one module: ps2, snes, and translator
